//////////////////////////////////////////////////////////////////////////////////
// Company: ITESO
// Engineer: Jorge Alberto Padilla Gutierrez
// Module Description: RISC-V ALU definitions
//////////////////////////////////////////////////////////////////////////////////

`define SEL_ADD     5'b00000
`define SEL_SUB	    5'b10000
`define SEL_XOR	    5'b00100
`define SEL_OR      5'b00110
`define SEL_AND	    5'b00111
`define SEL_SLL	    5'b00001
`define SEL_SRL	    5'b00101
`define SEL_SRA	    5'b10101
`define SEL_SLT	    5'b00010
`define SEL_SLTU	5'b00011
`define SEL_MUL     5'b01000